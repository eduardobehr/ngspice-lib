.title PWM with arbitrary non-linear source

.include pwm_generator.lib

* Generate input signals
Vfreq     freq        gnd       2000
Vsine     signal      gnd       SIN(0 1 60)

* Feed signals to pwm generator
xpwm      signal      freq      pwm          PWM3

* Filter output
.param order = 1

.if (order == 1)
  Rf        pwm         filtered  1000
  Cf        filtered    gnd       1u
.elseif (order == 2)
  Lf1       pwm         cap       1n
  Cf        cap         gnd       1u
  Lf2       cap         filtered  1n
.endif

.tran 1u 20m

.control
  run
  plot v(signal) v(pwm) filtered
.endc