.title Test SPDT
*
* This test circuit puts an inductor in series with the SPDT switch's terminal 1
*   in order to verify state continuity after switching. 
*

.include SPDT.lib
.include ../../diode/ideal/idiode.lib

** Command pulses generation
Vs      cmd     gnd     PULSE(0 2 2NS 2NS 2NS 80us 100us)

** Input stage
Vin     3       gnd     48

** Switch under test
Xsw     1       gnd     3       cmd     SPDT
  
** Output stage
L1      1       out     2000uH
RL      out     gnd     5
* Note: there is no need for a diode!


.tran 1us 100ms uic


.control
    run
    plot l1#branch
.endc
