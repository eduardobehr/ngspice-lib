PWM with arbitrary non-linear source

.param sawtooth_period = 0.0001


R1              vcc             gnd     10

BsawtoothP      sawtoothP       gnd     v=0.5+(time/sawtooth_period-floor(0.5+time/sawtooth_period))
BsawtoothM      sawtoothM       gnd     v=-0.5+(time/sawtooth_period-floor(0.5+time/sawtooth_period))
Binputsine      sine            gnd     v=sin(time*2*3.141593*60)
Bpwm            pwm             gnd     v=v(sine)>=v(sawtoothP) && v(sine)>=0 ? 1 : v(sine)<=v(sawtoothM) && v(sine)<=0 ? -1 : 0


.tran 1u 20m

.control
  run
  plot sine sawtoothP sawtoothM
  plot pwm
.endc