.title Test exp
.include exponentiation.lib

** Input signals
bV1      sig1    gnd     v={1*sin(377*time)}
V2      sig2    gnd     3

** Output signals
*
X_12   sig1   sig2   outvar      YEXPX_VAR
*
X_23   sig1   outfix      YEXPX_FIX x=2

.tran 1us 10m uic

.control
    run
    plot sig1 outvar outfix
.endc
