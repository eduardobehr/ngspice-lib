.title Test exp
.include exponentiation.lib

** Input signals
V1      sig1    gnd     -2
V2      sig2    gnd     3

** Output signals
*
X_12   sig1   sig2   out1      YEXPX_VAR
*
X_23   sig1   out2      YEXPX_FIX x=2

.tran

.control
    run
    plot sig1 out1 out2
.endc
